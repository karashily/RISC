library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;

entity RAM is
  port(
   RAM_CLOCK: in std_logic; 
   RAM_INS_ADDR: in std_logic_vector(10 downto 0);  
   RAM_DATA_ADDR: in std_logic_vector(10 downto 0);  
   RAM_DATA_WR: in std_logic;
   RAM_INS_WR: in std_logic; 
   RAM_INS_IN: in std_logic_vector(15 downto 0);
   RAM_INS_OUT: out std_logic_vector(15 downto 0);
   RAM_DATA_IN: in std_logic_vector(31 downto 0);
   RAM_DATA_OUT: out std_logic_vector(31 downto 0)
  );
end RAM;

architecture Behavioral of RAM is
type RAM_ARRAY is array (0 to 2047 ) of std_logic_vector (15 downto 0);
signal RAM: RAM_ARRAY :=(
  0 => "0000000000010000",
  1 => "0000000000000000",
  2 => "0000000100000000",
  3 => "0000000000000000",
  4 => "0100000000000000",
  5 => "0100000000000000",
  6 => "0100000000000000",
  7 => "0100000000000000",
  8 => "0100000000000000",
  9 => "0100000000000000",
  10 => "0100000000000000",
  11 => "0100000000000000",
  12 => "0100000000000000",
  13 => "0100000000000000",
  14 => "0100000000000000",
  15 => "0100000000000000",
  16 => "0110100100000000",
  17 => "0110101000000000",
  18 => "0110101100000000",
  19 => "0110110000000000",
  20 => "0110111000000000",
  21 => "0110111100000000",
  22 => "1000010000000000",
  23 => "1100100100000000",
  24 => "0101011100000000",
  25 => "0100000000000000",
  26 => "0100000000000000",
  27 => "0100000000000000",
  28 => "0100000000000000",
  29 => "0100000000000000",
  30 => "0100000000000000",
  31 => "0100000000000000",
  32 => "0100000000000000",
  33 => "0100000000000000",
  34 => "0100000000000000",
  35 => "0100000000000000",
  36 => "0100000000000000",
  37 => "0100000000000000",
  38 => "0100000000000000",
  39 => "0100000000000000",
  40 => "0100000000000000",
  41 => "0100000000000000",
  42 => "0100000000000000",
  43 => "0100000000000000",
  44 => "0100000000000000",
  45 => "0100000000000000",
  46 => "0100000000000000",
  47 => "0100000000000000",
  48 => "0001100110110100",
  49 => "1100001000000000",
  50 => "0101011100000000",
  51 => "0100000000000000",
  52 => "0100000000000000",
  53 => "0100000000000000",
  54 => "0100000000000000",
  55 => "0100000000000000",
  56 => "0100000000000000",
  57 => "0100000000000000",
  58 => "0100000000000000",
  59 => "0100000000000000",
  60 => "0100000000000000",
  61 => "0100000000000000",
  62 => "0100000000000000",
  63 => "0100000000000000",
  64 => "0100000000000000",
  65 => "0100000000000000",
  66 => "0100000000000000",
  67 => "0100000000000000",
  68 => "0100000000000000",
  69 => "0100000000000000",
  70 => "0100000000000000",
  71 => "0100000000000000",
  72 => "0100000000000000",
  73 => "0100000000000000",
  74 => "0100000000000000",
  75 => "0100000000000000",
  76 => "0100000000000000",
  77 => "0100000000000000",
  78 => "0100000000000000",
  79 => "0100000000000000",
  80 => "1100001100000000",
  81 => "0100110100000000",
  82 => "0101010100000000",
  83 => "0110111000000000",
  84 => "1100011000000000",
  85 => "0101000100000000",
  86 => "0100000000000000",
  87 => "0100000000000000",
  88 => "0100000000000000",
  89 => "0100000000000000",
  90 => "0100000000000000",
  91 => "0100000000000000",
  92 => "0100000000000000",
  93 => "0100000000000000",
  94 => "0100000000000000",
  95 => "0100000000000000",
  96 => "0100000000000000",
  97 => "0100000000000000",
  98 => "0100000000000000",
  99 => "0100000000000000",
  100 => "0100000000000000",
  101 => "0100000000000000",
  102 => "0100000000000000",
  103 => "0100000000000000",
  104 => "0100000000000000",
  105 => "0100000000000000",
  106 => "0100000000000000",
  107 => "0100000000000000",
  108 => "0100000000000000",
  109 => "0100000000000000",
  110 => "0100000000000000",
  111 => "0100000000000000",
  112 => "0100000000000000",
  113 => "0100000000000000",
  114 => "0100000000000000",
  115 => "0100000000000000",
  116 => "0100000000000000",
  117 => "0100000000000000",
  118 => "0100000000000000",
  119 => "0100000000000000",
  120 => "0100000000000000",
  121 => "0100000000000000",
  122 => "0100000000000000",
  123 => "0100000000000000",
  124 => "0100000000000000",
  125 => "0100000000000000",
  126 => "0100000000000000",
  127 => "0100000000000000",
  128 => "0100000000000000",
  129 => "0100000000000000",
  130 => "0100000000000000",
  131 => "0100000000000000",
  132 => "0100000000000000",
  133 => "0100000000000000",
  134 => "0100000000000000",
  135 => "0100000000000000",
  136 => "0100000000000000",
  137 => "0100000000000000",
  138 => "0100000000000000",
  139 => "0100000000000000",
  140 => "0100000000000000",
  141 => "0100000000000000",
  142 => "0100000000000000",
  143 => "0100000000000000",
  144 => "0100000000000000",
  145 => "0100000000000000",
  146 => "0100000000000000",
  147 => "0100000000000000",
  148 => "0100000000000000",
  149 => "0100000000000000",
  150 => "0100000000000000",
  151 => "0100000000000000",
  152 => "0100000000000000",
  153 => "0100000000000000",
  154 => "0100000000000000",
  155 => "0100000000000000",
  156 => "0100000000000000",
  157 => "0100000000000000",
  158 => "0100000000000000",
  159 => "0100000000000000",
  160 => "0100000000000000",
  161 => "0100000000000000",
  162 => "0100000000000000",
  163 => "0100000000000000",
  164 => "0100000000000000",
  165 => "0100000000000000",
  166 => "0100000000000000",
  167 => "0100000000000000",
  168 => "0100000000000000",
  169 => "0100000000000000",
  170 => "0100000000000000",
  171 => "0100000000000000",
  172 => "0100000000000000",
  173 => "0100000000000000",
  174 => "0100000000000000",
  175 => "0100000000000000",
  176 => "0100000000000000",
  177 => "0100000000000000",
  178 => "0100000000000000",
  179 => "0100000000000000",
  180 => "0100000000000000",
  181 => "0100000000000000",
  182 => "0100000000000000",
  183 => "0100000000000000",
  184 => "0100000000000000",
  185 => "0100000000000000",
  186 => "0100000000000000",
  187 => "0100000000000000",
  188 => "0100000000000000",
  189 => "0100000000000000",
  190 => "0100000000000000",
  191 => "0100000000000000",
  192 => "0100000000000000",
  193 => "0100000000000000",
  194 => "0100000000000000",
  195 => "0100000000000000",
  196 => "0100000000000000",
  197 => "0100000000000000",
  198 => "0100000000000000",
  199 => "0100000000000000",
  200 => "0100000000000000",
  201 => "0100000000000000",
  202 => "0100000000000000",
  203 => "0100000000000000",
  204 => "0100000000000000",
  205 => "0100000000000000",
  206 => "0100000000000000",
  207 => "0100000000000000",
  208 => "0100000000000000",
  209 => "0100000000000000",
  210 => "0100000000000000",
  211 => "0100000000000000",
  212 => "0100000000000000",
  213 => "0100000000000000",
  214 => "0100000000000000",
  215 => "0100000000000000",
  216 => "0100000000000000",
  217 => "0100000000000000",
  218 => "0100000000000000",
  219 => "0100000000000000",
  220 => "0100000000000000",
  221 => "0100000000000000",
  222 => "0100000000000000",
  223 => "0100000000000000",
  224 => "0100000000000000",
  225 => "0100000000000000",
  226 => "0100000000000000",
  227 => "0100000000000000",
  228 => "0100000000000000",
  229 => "0100000000000000",
  230 => "0100000000000000",
  231 => "0100000000000000",
  232 => "0100000000000000",
  233 => "0100000000000000",
  234 => "0100000000000000",
  235 => "0100000000000000",
  236 => "0100000000000000",
  237 => "0100000000000000",
  238 => "0100000000000000",
  239 => "0100000000000000",
  240 => "0100000000000000",
  241 => "0100000000000000",
  242 => "0100000000000000",
  243 => "0100000000000000",
  244 => "0100000000000000",
  245 => "0100000000000000",
  246 => "0100000000000000",
  247 => "0100000000000000",
  248 => "0100000000000000",
  249 => "0100000000000000",
  250 => "0100000000000000",
  251 => "0100000000000000",
  252 => "0100000000000000",
  253 => "0100000000000000",
  254 => "0100000000000000",
  255 => "0100000000000000",
  256 => "0000000000000000",
  257 => "0110011000000000",
  258 => "1110000000000000",
  259 => "0100000000000000",
  260 => "0100000000000000",
  261 => "0100000000000000",
  262 => "0100000000000000",
  263 => "0100000000000000",
  264 => "0100000000000000",
  265 => "0100000000000000",
  266 => "0100000000000000",
  267 => "0100000000000000",
  268 => "0100000000000000",
  269 => "0100000000000000",
  270 => "0100000000000000",
  271 => "0100000000000000",
  272 => "0100000000000000",
  273 => "0100000000000000",
  274 => "0100000000000000",
  275 => "0100000000000000",
  276 => "0100000000000000",
  277 => "0100000000000000",
  278 => "0100000000000000",
  279 => "0100000000000000",
  280 => "0100000000000000",
  281 => "0100000000000000",
  282 => "0100000000000000",
  283 => "0100000000000000",
  284 => "0100000000000000",
  285 => "0100000000000000",
  286 => "0100000000000000",
  287 => "0100000000000000",
  288 => "0100000000000000",
  289 => "0100000000000000",
  290 => "0100000000000000",
  291 => "0100000000000000",
  292 => "0100000000000000",
  293 => "0100000000000000",
  294 => "0100000000000000",
  295 => "0100000000000000",
  296 => "0100000000000000",
  297 => "0100000000000000",
  298 => "0100000000000000",
  299 => "0100000000000000",
  300 => "0100000000000000",
  301 => "0100000000000000",
  302 => "0100000000000000",
  303 => "0100000000000000",
  304 => "0100000000000000",
  305 => "0100000000000000",
  306 => "0100000000000000",
  307 => "0100000000000000",
  308 => "0100000000000000",
  309 => "0100000000000000",
  310 => "0100000000000000",
  311 => "0100000000000000",
  312 => "0100000000000000",
  313 => "0100000000000000",
  314 => "0100000000000000",
  315 => "0100000000000000",
  316 => "0100000000000000",
  317 => "0100000000000000",
  318 => "0100000000000000",
  319 => "0100000000000000",
  320 => "0100000000000000",
  321 => "0100000000000000",
  322 => "0100000000000000",
  323 => "0100000000000000",
  324 => "0100000000000000",
  325 => "0100000000000000",
  326 => "0100000000000000",
  327 => "0100000000000000",
  328 => "0100000000000000",
  329 => "0100000000000000",
  330 => "0100000000000000",
  331 => "0100000000000000",
  332 => "0100000000000000",
  333 => "0100000000000000",
  334 => "0100000000000000",
  335 => "0100000000000000",
  336 => "0100000000000000",
  337 => "0100000000000000",
  338 => "0100000000000000",
  339 => "0100000000000000",
  340 => "0100000000000000",
  341 => "0100000000000000",
  342 => "0100000000000000",
  343 => "0100000000000000",
  344 => "0100000000000000",
  345 => "0100000000000000",
  346 => "0100000000000000",
  347 => "0100000000000000",
  348 => "0100000000000000",
  349 => "0100000000000000",
  350 => "0100000000000000",
  351 => "0100000000000000",
  352 => "0100000000000000",
  353 => "0100000000000000",
  354 => "0100000000000000",
  355 => "0100000000000000",
  356 => "0100000000000000",
  357 => "0100000000000000",
  358 => "0100000000000000",
  359 => "0100000000000000",
  360 => "0100000000000000",
  361 => "0100000000000000",
  362 => "0100000000000000",
  363 => "0100000000000000",
  364 => "0100000000000000",
  365 => "0100000000000000",
  366 => "0100000000000000",
  367 => "0100000000000000",
  368 => "0100000000000000",
  369 => "0100000000000000",
  370 => "0100000000000000",
  371 => "0100000000000000",
  372 => "0100000000000000",
  373 => "0100000000000000",
  374 => "0100000000000000",
  375 => "0100000000000000",
  376 => "0100000000000000",
  377 => "0100000000000000",
  378 => "0100000000000000",
  379 => "0100000000000000",
  380 => "0100000000000000",
  381 => "0100000000000000",
  382 => "0100000000000000",
  383 => "0100000000000000",
  384 => "0100000000000000",
  385 => "0100000000000000",
  386 => "0100000000000000",
  387 => "0100000000000000",
  388 => "0100000000000000",
  389 => "0100000000000000",
  390 => "0100000000000000",
  391 => "0100000000000000",
  392 => "0100000000000000",
  393 => "0100000000000000",
  394 => "0100000000000000",
  395 => "0100000000000000",
  396 => "0100000000000000",
  397 => "0100000000000000",
  398 => "0100000000000000",
  399 => "0100000000000000",
  400 => "0100000000000000",
  401 => "0100000000000000",
  402 => "0100000000000000",
  403 => "0100000000000000",
  404 => "0100000000000000",
  405 => "0100000000000000",
  406 => "0100000000000000",
  407 => "0100000000000000",
  408 => "0100000000000000",
  409 => "0100000000000000",
  410 => "0100000000000000",
  411 => "0100000000000000",
  412 => "0100000000000000",
  413 => "0100000000000000",
  414 => "0100000000000000",
  415 => "0100000000000000",
  416 => "0100000000000000",
  417 => "0100000000000000",
  418 => "0100000000000000",
  419 => "0100000000000000",
  420 => "0100000000000000",
  421 => "0100000000000000",
  422 => "0100000000000000",
  423 => "0100000000000000",
  424 => "0100000000000000",
  425 => "0100000000000000",
  426 => "0100000000000000",
  427 => "0100000000000000",
  428 => "0100000000000000",
  429 => "0100000000000000",
  430 => "0100000000000000",
  431 => "0100000000000000",
  432 => "0100000000000000",
  433 => "0100000000000000",
  434 => "0100000000000000",
  435 => "0100000000000000",
  436 => "0100000000000000",
  437 => "0100000000000000",
  438 => "0100000000000000",
  439 => "0100000000000000",
  440 => "0100000000000000",
  441 => "0100000000000000",
  442 => "0100000000000000",
  443 => "0100000000000000",
  444 => "0100000000000000",
  445 => "0100000000000000",
  446 => "0100000000000000",
  447 => "0100000000000000",
  448 => "0100000000000000",
  449 => "0100000000000000",
  450 => "0100000000000000",
  451 => "0100000000000000",
  452 => "0100000000000000",
  453 => "0100000000000000",
  454 => "0100000000000000",
  455 => "0100000000000000",
  456 => "0100000000000000",
  457 => "0100000000000000",
  458 => "0100000000000000",
  459 => "0100000000000000",
  460 => "0100000000000000",
  461 => "0100000000000000",
  462 => "0100000000000000",
  463 => "0100000000000000",
  464 => "0100000000000000",
  465 => "0100000000000000",
  466 => "0100000000000000",
  467 => "0100000000000000",
  468 => "0100000000000000",
  469 => "0100000000000000",
  470 => "0100000000000000",
  471 => "0100000000000000",
  472 => "0100000000000000",
  473 => "0100000000000000",
  474 => "0100000000000000",
  475 => "0100000000000000",
  476 => "0100000000000000",
  477 => "0100000000000000",
  478 => "0100000000000000",
  479 => "0100000000000000",
  480 => "0100000000000000",
  481 => "0100000000000000",
  482 => "0100000000000000",
  483 => "0100000000000000",
  484 => "0100000000000000",
  485 => "0100000000000000",
  486 => "0100000000000000",
  487 => "0100000000000000",
  488 => "0100000000000000",
  489 => "0100000000000000",
  490 => "0100000000000000",
  491 => "0100000000000000",
  492 => "0100000000000000",
  493 => "0100000000000000",
  494 => "0100000000000000",
  495 => "0100000000000000",
  496 => "0100000000000000",
  497 => "0100000000000000",
  498 => "0100000000000000",
  499 => "0100000000000000",
  500 => "0100000000000000",
  501 => "0100000000000000",
  502 => "0100000000000000",
  503 => "0100000000000000",
  504 => "0100000000000000",
  505 => "0100000000000000",
  506 => "0100000000000000",
  507 => "0100000000000000",
  508 => "0100000000000000",
  509 => "0100000000000000",
  510 => "0100000000000000",
  511 => "0100000000000000",
  512 => "1000111000000000",
  513 => "1101011000000000",
  514 => "0101011000000000",
  515 => "0100000000000000",
  516 => "0100000000000000",
  517 => "0100000000000000",
  518 => "0100000000000000",
  519 => "0100000000000000",
  520 => "0100000000000000",
  521 => "0100000000000000",
  522 => "0100000000000000",
  523 => "0100000000000000",
  524 => "0100000000000000",
  525 => "0100000000000000",
  526 => "0100000000000000",
  527 => "0100000000000000",
  528 => "0100000000000000",
  529 => "0100000000000000",
  530 => "0100000000000000",
  531 => "0100000000000000",
  532 => "0100000000000000",
  533 => "0100000000000000",
  534 => "0100000000000000",
  535 => "0100000000000000",
  536 => "0100000000000000",
  537 => "0100000000000000",
  538 => "0100000000000000",
  539 => "0100000000000000",
  540 => "0100000000000000",
  541 => "0100000000000000",
  542 => "0100000000000000",
  543 => "0100000000000000",
  544 => "0100000000000000",
  545 => "0100000000000000",
  546 => "0100000000000000",
  547 => "0100000000000000",
  548 => "0100000000000000",
  549 => "0100000000000000",
  550 => "0100000000000000",
  551 => "0100000000000000",
  552 => "0100000000000000",
  553 => "0100000000000000",
  554 => "0100000000000000",
  555 => "0100000000000000",
  556 => "0100000000000000",
  557 => "0100000000000000",
  558 => "0100000000000000",
  559 => "0100000000000000",
  560 => "0100000000000000",
  561 => "0100000000000000",
  562 => "0100000000000000",
  563 => "0100000000000000",
  564 => "0100000000000000",
  565 => "0100000000000000",
  566 => "0100000000000000",
  567 => "0100000000000000",
  568 => "0100000000000000",
  569 => "0100000000000000",
  570 => "0100000000000000",
  571 => "0100000000000000",
  572 => "0100000000000000",
  573 => "0100000000000000",
  574 => "0100000000000000",
  575 => "0100000000000000",
  576 => "0100000000000000",
  577 => "0100000000000000",
  578 => "0100000000000000",
  579 => "0100000000000000",
  580 => "0100000000000000",
  581 => "0100000000000000",
  582 => "0100000000000000",
  583 => "0100000000000000",
  584 => "0100000000000000",
  585 => "0100000000000000",
  586 => "0100000000000000",
  587 => "0100000000000000",
  588 => "0100000000000000",
  589 => "0100000000000000",
  590 => "0100000000000000",
  591 => "0100000000000000",
  592 => "0100000000000000",
  593 => "0100000000000000",
  594 => "0100000000000000",
  595 => "0100000000000000",
  596 => "0100000000000000",
  597 => "0100000000000000",
  598 => "0100000000000000",
  599 => "0100000000000000",
  600 => "0100000000000000",
  601 => "0100000000000000",
  602 => "0100000000000000",
  603 => "0100000000000000",
  604 => "0100000000000000",
  605 => "0100000000000000",
  606 => "0100000000000000",
  607 => "0100000000000000",
  608 => "0100000000000000",
  609 => "0100000000000000",
  610 => "0100000000000000",
  611 => "0100000000000000",
  612 => "0100000000000000",
  613 => "0100000000000000",
  614 => "0100000000000000",
  615 => "0100000000000000",
  616 => "0100000000000000",
  617 => "0100000000000000",
  618 => "0100000000000000",
  619 => "0100000000000000",
  620 => "0100000000000000",
  621 => "0100000000000000",
  622 => "0100000000000000",
  623 => "0100000000000000",
  624 => "0100000000000000",
  625 => "0100000000000000",
  626 => "0100000000000000",
  627 => "0100000000000000",
  628 => "0100000000000000",
  629 => "0100000000000000",
  630 => "0100000000000000",
  631 => "0100000000000000",
  632 => "0100000000000000",
  633 => "0100000000000000",
  634 => "0100000000000000",
  635 => "0100000000000000",
  636 => "0100000000000000",
  637 => "0100000000000000",
  638 => "0100000000000000",
  639 => "0100000000000000",
  640 => "0100000000000000",
  641 => "0100000000000000",
  642 => "0100000000000000",
  643 => "0100000000000000",
  644 => "0100000000000000",
  645 => "0100000000000000",
  646 => "0100000000000000",
  647 => "0100000000000000",
  648 => "0100000000000000",
  649 => "0100000000000000",
  650 => "0100000000000000",
  651 => "0100000000000000",
  652 => "0100000000000000",
  653 => "0100000000000000",
  654 => "0100000000000000",
  655 => "0100000000000000",
  656 => "0100000000000000",
  657 => "0100000000000000",
  658 => "0100000000000000",
  659 => "0100000000000000",
  660 => "0100000000000000",
  661 => "0100000000000000",
  662 => "0100000000000000",
  663 => "0100000000000000",
  664 => "0100000000000000",
  665 => "0100000000000000",
  666 => "0100000000000000",
  667 => "0100000000000000",
  668 => "0100000000000000",
  669 => "0100000000000000",
  670 => "0100000000000000",
  671 => "0100000000000000",
  672 => "0100000000000000",
  673 => "0100000000000000",
  674 => "0100000000000000",
  675 => "0100000000000000",
  676 => "0100000000000000",
  677 => "0100000000000000",
  678 => "0100000000000000",
  679 => "0100000000000000",
  680 => "0100000000000000",
  681 => "0100000000000000",
  682 => "0100000000000000",
  683 => "0100000000000000",
  684 => "0100000000000000",
  685 => "0100000000000000",
  686 => "0100000000000000",
  687 => "0100000000000000",
  688 => "0100000000000000",
  689 => "0100000000000000",
  690 => "0100000000000000",
  691 => "0100000000000000",
  692 => "0100000000000000",
  693 => "0100000000000000",
  694 => "0100000000000000",
  695 => "0100000000000000",
  696 => "0100000000000000",
  697 => "0100000000000000",
  698 => "0100000000000000",
  699 => "0100000000000000",
  700 => "0100000000000000",
  701 => "0100000000000000",
  702 => "0100000000000000",
  703 => "0100000000000000",
  704 => "0100000000000000",
  705 => "0100000000000000",
  706 => "0100000000000000",
  707 => "0100000000000000",
  708 => "0100000000000000",
  709 => "0100000000000000",
  710 => "0100000000000000",
  711 => "0100000000000000",
  712 => "0100000000000000",
  713 => "0100000000000000",
  714 => "0100000000000000",
  715 => "0100000000000000",
  716 => "0100000000000000",
  717 => "0100000000000000",
  718 => "0100000000000000",
  719 => "0100000000000000",
  720 => "0100000000000000",
  721 => "0100000000000000",
  722 => "0100000000000000",
  723 => "0100000000000000",
  724 => "0100000000000000",
  725 => "0100000000000000",
  726 => "0100000000000000",
  727 => "0100000000000000",
  728 => "0100000000000000",
  729 => "0100000000000000",
  730 => "0100000000000000",
  731 => "0100000000000000",
  732 => "0100000000000000",
  733 => "0100000000000000",
  734 => "0100000000000000",
  735 => "0100000000000000",
  736 => "0100000000000000",
  737 => "0100000000000000",
  738 => "0100000000000000",
  739 => "0100000000000000",
  740 => "0100000000000000",
  741 => "0100000000000000",
  742 => "0100000000000000",
  743 => "0100000000000000",
  744 => "0100000000000000",
  745 => "0100000000000000",
  746 => "0100000000000000",
  747 => "0100000000000000",
  748 => "0100000000000000",
  749 => "0100000000000000",
  750 => "0100000000000000",
  751 => "0100000000000000",
  752 => "0100000000000000",
  753 => "0100000000000000",
  754 => "0100000000000000",
  755 => "0100000000000000",
  756 => "0100000000000000",
  757 => "0100000000000000",
  758 => "0100000000000000",
  759 => "0100000000000000",
  760 => "0100000000000000",
  761 => "0100000000000000",
  762 => "0100000000000000",
  763 => "0100000000000000",
  764 => "0100000000000000",
  765 => "0100000000000000",
  766 => "0100000000000000",
  767 => "0100000000000000",
  768 => "0000001111011000",
  769 => "0000000101000100",
  770 => "1101100000000000",
  771 => "0101011100000000",
  772 => "0100000000000000",
  773 => "0100000000000000",
  774 => "0100000000000000",
  775 => "0100000000000000",
  776 => "0100000000000000",
  777 => "0100000000000000",
  778 => "0100000000000000",
  779 => "0100000000000000",
  780 => "0100000000000000",
  781 => "0100000000000000",
  782 => "0100000000000000",
  783 => "0100000000000000",
  784 => "0100000000000000",
  785 => "0100000000000000",
  786 => "0100000000000000",
  787 => "0100000000000000",
  788 => "0100000000000000",
  789 => "0100000000000000",
  790 => "0100000000000000",
  791 => "0100000000000000",
  792 => "0100000000000000",
  793 => "0100000000000000",
  794 => "0100000000000000",
  795 => "0100000000000000",
  796 => "0100000000000000",
  797 => "0100000000000000",
  798 => "0100000000000000",
  799 => "0100000000000000",
  800 => "0100000000000000",
  801 => "0100000000000000",
  802 => "0100000000000000",
  803 => "0100000000000000",
  804 => "0100000000000000",
  805 => "0100000000000000",
  806 => "0100000000000000",
  807 => "0100000000000000",
  808 => "0100000000000000",
  809 => "0100000000000000",
  810 => "0100000000000000",
  811 => "0100000000000000",
  812 => "0100000000000000",
  813 => "0100000000000000",
  814 => "0100000000000000",
  815 => "0100000000000000",
  816 => "0100000000000000",
  817 => "0100000000000000",
  818 => "0100000000000000",
  819 => "0100000000000000",
  820 => "0100000000000000",
  821 => "0100000000000000",
  822 => "0100000000000000",
  823 => "0100000000000000",
  824 => "0100000000000000",
  825 => "0100000000000000",
  826 => "0100000000000000",
  827 => "0100000000000000",
  828 => "0100000000000000",
  829 => "0100000000000000",
  830 => "0100000000000000",
  831 => "0100000000000000",
  832 => "0100000000000000",
  833 => "0100000000000000",
  834 => "0100000000000000",
  835 => "0100000000000000",
  836 => "0100000000000000",
  837 => "0100000000000000",
  838 => "0100000000000000",
  839 => "0100000000000000",
  840 => "0100000000000000",
  841 => "0100000000000000",
  842 => "0100000000000000",
  843 => "0100000000000000",
  844 => "0100000000000000",
  845 => "0100000000000000",
  846 => "0100000000000000",
  847 => "0100000000000000",
  848 => "0100000000000000",
  849 => "0100000000000000",
  850 => "0100000000000000",
  851 => "0100000000000000",
  852 => "0100000000000000",
  853 => "0100000000000000",
  854 => "0100000000000000",
  855 => "0100000000000000",
  856 => "0100000000000000",
  857 => "0100000000000000",
  858 => "0100000000000000",
  859 => "0100000000000000",
  860 => "0100000000000000",
  861 => "0100000000000000",
  862 => "0100000000000000",
  863 => "0100000000000000",
  864 => "0100000000000000",
  865 => "0100000000000000",
  866 => "0100000000000000",
  867 => "0100000000000000",
  868 => "0100000000000000",
  869 => "0100000000000000",
  870 => "0100000000000000",
  871 => "0100000000000000",
  872 => "0100000000000000",
  873 => "0100000000000000",
  874 => "0100000000000000",
  875 => "0100000000000000",
  876 => "0100000000000000",
  877 => "0100000000000000",
  878 => "0100000000000000",
  879 => "0100000000000000",
  880 => "0100000000000000",
  881 => "0100000000000000",
  882 => "0100000000000000",
  883 => "0100000000000000",
  884 => "0100000000000000",
  885 => "0100000000000000",
  886 => "0100000000000000",
  887 => "0100000000000000",
  888 => "0100000000000000",
  889 => "0100000000000000",
  890 => "0100000000000000",
  891 => "0100000000000000",
  892 => "0100000000000000",
  893 => "0100000000000000",
  894 => "0100000000000000",
  895 => "0100000000000000",
  896 => "0100000000000000",
  897 => "0100000000000000",
  898 => "0100000000000000",
  899 => "0100000000000000",
  900 => "0100000000000000",
  901 => "0100000000000000",
  902 => "0100000000000000",
  903 => "0100000000000000",
  904 => "0100000000000000",
  905 => "0100000000000000",
  906 => "0100000000000000",
  907 => "0100000000000000",
  908 => "0100000000000000",
  909 => "0100000000000000",
  910 => "0100000000000000",
  911 => "0100000000000000",
  912 => "0100000000000000",
  913 => "0100000000000000",
  914 => "0100000000000000",
  915 => "0100000000000000",
  916 => "0100000000000000",
  917 => "0100000000000000",
  918 => "0100000000000000",
  919 => "0100000000000000",
  920 => "0100000000000000",
  921 => "0100000000000000",
  922 => "0100000000000000",
  923 => "0100000000000000",
  924 => "0100000000000000",
  925 => "0100000000000000",
  926 => "0100000000000000",
  927 => "0100000000000000",
  928 => "0100000000000000",
  929 => "0100000000000000",
  930 => "0100000000000000",
  931 => "0100000000000000",
  932 => "0100000000000000",
  933 => "0100000000000000",
  934 => "0100000000000000",
  935 => "0100000000000000",
  936 => "0100000000000000",
  937 => "0100000000000000",
  938 => "0100000000000000",
  939 => "0100000000000000",
  940 => "0100000000000000",
  941 => "0100000000000000",
  942 => "0100000000000000",
  943 => "0100000000000000",
  944 => "0100000000000000",
  945 => "0100000000000000",
  946 => "0100000000000000",
  947 => "0100000000000000",
  948 => "0100000000000000",
  949 => "0100000000000000",
  950 => "0100000000000000",
  951 => "0100000000000000",
  952 => "0100000000000000",
  953 => "0100000000000000",
  954 => "0100000000000000",
  955 => "0100000000000000",
  956 => "0100000000000000",
  957 => "0100000000000000",
  958 => "0100000000000000",
  959 => "0100000000000000",
  960 => "0100000000000000",
  961 => "0100000000000000",
  962 => "0100000000000000",
  963 => "0100000000000000",
  964 => "0100000000000000",
  965 => "0100000000000000",
  966 => "0100000000000000",
  967 => "0100000000000000",
  968 => "0100000000000000",
  969 => "0100000000000000",
  970 => "0100000000000000",
  971 => "0100000000000000",
  972 => "0100000000000000",
  973 => "0100000000000000",
  974 => "0100000000000000",
  975 => "0100000000000000",
  976 => "0100000000000000",
  977 => "0100000000000000",
  978 => "0100000000000000",
  979 => "0100000000000000",
  980 => "0100000000000000",
  981 => "0100000000000000",
  982 => "0100000000000000",
  983 => "0100000000000000",
  984 => "0100000000000000",
  985 => "0100000000000000",
  986 => "0100000000000000",
  987 => "0100000000000000",
  988 => "0100000000000000",
  989 => "0100000000000000",
  990 => "0100000000000000",
  991 => "0100000000000000",
  992 => "0100000000000000",
  993 => "0100000000000000",
  994 => "0100000000000000",
  995 => "0100000000000000",
  996 => "0100000000000000",
  997 => "0100000000000000",
  998 => "0100000000000000",
  999 => "0100000000000000",
  1000 => "0100000000000000",
  1001 => "0100000000000000",
  1002 => "0100000000000000",
  1003 => "0100000000000000",
  1004 => "0100000000000000",
  1005 => "0100000000000000",
  1006 => "0100000000000000",
  1007 => "0100000000000000",
  1008 => "0100000000000000",
  1009 => "0100000000000000",
  1010 => "0100000000000000",
  1011 => "0100000000000000",
  1012 => "0100000000000000",
  1013 => "0100000000000000",
  1014 => "0100000000000000",
  1015 => "0100000000000000",
  1016 => "0100000000000000",
  1017 => "0100000000000000",
  1018 => "0100000000000000",
  1019 => "0100000000000000",
  1020 => "0100000000000000",
  1021 => "0100000000000000",
  1022 => "0100000000000000",
  1023 => "0100000000000000",
  1024 => "0100000000000000",
  1025 => "0100000000000000",
  1026 => "0100000000000000",
  1027 => "0100000000000000",
  1028 => "0100000000000000",
  1029 => "0100000000000000",
  1030 => "0100000000000000",
  1031 => "0100000000000000",
  1032 => "0100000000000000",
  1033 => "0100000000000000",
  1034 => "0100000000000000",
  1035 => "0100000000000000",
  1036 => "0100000000000000",
  1037 => "0100000000000000",
  1038 => "0100000000000000",
  1039 => "0100000000000000",
  1040 => "0100000000000000",
  1041 => "0100000000000000",
  1042 => "0100000000000000",
  1043 => "0100000000000000",
  1044 => "0100000000000000",
  1045 => "0100000000000000",
  1046 => "0100000000000000",
  1047 => "0100000000000000",
  1048 => "0100000000000000",
  1049 => "0100000000000000",
  1050 => "0100000000000000",
  1051 => "0100000000000000",
  1052 => "0100000000000000",
  1053 => "0100000000000000",
  1054 => "0100000000000000",
  1055 => "0100000000000000",
  1056 => "0100000000000000",
  1057 => "0100000000000000",
  1058 => "0100000000000000",
  1059 => "0100000000000000",
  1060 => "0100000000000000",
  1061 => "0100000000000000",
  1062 => "0100000000000000",
  1063 => "0100000000000000",
  1064 => "0100000000000000",
  1065 => "0100000000000000",
  1066 => "0100000000000000",
  1067 => "0100000000000000",
  1068 => "0100000000000000",
  1069 => "0100000000000000",
  1070 => "0100000000000000",
  1071 => "0100000000000000",
  1072 => "0100000000000000",
  1073 => "0100000000000000",
  1074 => "0100000000000000",
  1075 => "0100000000000000",
  1076 => "0100000000000000",
  1077 => "0100000000000000",
  1078 => "0100000000000000",
  1079 => "0100000000000000",
  1080 => "0100000000000000",
  1081 => "0100000000000000",
  1082 => "0100000000000000",
  1083 => "0100000000000000",
  1084 => "0100000000000000",
  1085 => "0100000000000000",
  1086 => "0100000000000000",
  1087 => "0100000000000000",
  1088 => "0100000000000000",
  1089 => "0100000000000000",
  1090 => "0100000000000000",
  1091 => "0100000000000000",
  1092 => "0100000000000000",
  1093 => "0100000000000000",
  1094 => "0100000000000000",
  1095 => "0100000000000000",
  1096 => "0100000000000000",
  1097 => "0100000000000000",
  1098 => "0100000000000000",
  1099 => "0100000000000000",
  1100 => "0100000000000000",
  1101 => "0100000000000000",
  1102 => "0100000000000000",
  1103 => "0100000000000000",
  1104 => "0100000000000000",
  1105 => "0100000000000000",
  1106 => "0100000000000000",
  1107 => "0100000000000000",
  1108 => "0100000000000000",
  1109 => "0100000000000000",
  1110 => "0100000000000000",
  1111 => "0100000000000000",
  1112 => "0100000000000000",
  1113 => "0100000000000000",
  1114 => "0100000000000000",
  1115 => "0100000000000000",
  1116 => "0100000000000000",
  1117 => "0100000000000000",
  1118 => "0100000000000000",
  1119 => "0100000000000000",
  1120 => "0100000000000000",
  1121 => "0100000000000000",
  1122 => "0100000000000000",
  1123 => "0100000000000000",
  1124 => "0100000000000000",
  1125 => "0100000000000000",
  1126 => "0100000000000000",
  1127 => "0100000000000000",
  1128 => "0100000000000000",
  1129 => "0100000000000000",
  1130 => "0100000000000000",
  1131 => "0100000000000000",
  1132 => "0100000000000000",
  1133 => "0100000000000000",
  1134 => "0100000000000000",
  1135 => "0100000000000000",
  1136 => "0100000000000000",
  1137 => "0100000000000000",
  1138 => "0100000000000000",
  1139 => "0100000000000000",
  1140 => "0100000000000000",
  1141 => "0100000000000000",
  1142 => "0100000000000000",
  1143 => "0100000000000000",
  1144 => "0100000000000000",
  1145 => "0100000000000000",
  1146 => "0100000000000000",
  1147 => "0100000000000000",
  1148 => "0100000000000000",
  1149 => "0100000000000000",
  1150 => "0100000000000000",
  1151 => "0100000000000000",
  1152 => "0100000000000000",
  1153 => "0100000000000000",
  1154 => "0100000000000000",
  1155 => "0100000000000000",
  1156 => "0100000000000000",
  1157 => "0100000000000000",
  1158 => "0100000000000000",
  1159 => "0100000000000000",
  1160 => "0100000000000000",
  1161 => "0100000000000000",
  1162 => "0100000000000000",
  1163 => "0100000000000000",
  1164 => "0100000000000000",
  1165 => "0100000000000000",
  1166 => "0100000000000000",
  1167 => "0100000000000000",
  1168 => "0100000000000000",
  1169 => "0100000000000000",
  1170 => "0100000000000000",
  1171 => "0100000000000000",
  1172 => "0100000000000000",
  1173 => "0100000000000000",
  1174 => "0100000000000000",
  1175 => "0100000000000000",
  1176 => "0100000000000000",
  1177 => "0100000000000000",
  1178 => "0100000000000000",
  1179 => "0100000000000000",
  1180 => "0100000000000000",
  1181 => "0100000000000000",
  1182 => "0100000000000000",
  1183 => "0100000000000000",
  1184 => "0100000000000000",
  1185 => "0100000000000000",
  1186 => "0100000000000000",
  1187 => "0100000000000000",
  1188 => "0100000000000000",
  1189 => "0100000000000000",
  1190 => "0100000000000000",
  1191 => "0100000000000000",
  1192 => "0100000000000000",
  1193 => "0100000000000000",
  1194 => "0100000000000000",
  1195 => "0100000000000000",
  1196 => "0100000000000000",
  1197 => "0100000000000000",
  1198 => "0100000000000000",
  1199 => "0100000000000000",
  1200 => "0100000000000000",
  1201 => "0100000000000000",
  1202 => "0100000000000000",
  1203 => "0100000000000000",
  1204 => "0100000000000000",
  1205 => "0100000000000000",
  1206 => "0100000000000000",
  1207 => "0100000000000000",
  1208 => "0100000000000000",
  1209 => "0100000000000000",
  1210 => "0100000000000000",
  1211 => "0100000000000000",
  1212 => "0100000000000000",
  1213 => "0100000000000000",
  1214 => "0100000000000000",
  1215 => "0100000000000000",
  1216 => "0100000000000000",
  1217 => "0100000000000000",
  1218 => "0100000000000000",
  1219 => "0100000000000000",
  1220 => "0100000000000000",
  1221 => "0100000000000000",
  1222 => "0100000000000000",
  1223 => "0100000000000000",
  1224 => "0100000000000000",
  1225 => "0100000000000000",
  1226 => "0100000000000000",
  1227 => "0100000000000000",
  1228 => "0100000000000000",
  1229 => "0100000000000000",
  1230 => "0100000000000000",
  1231 => "0100000000000000",
  1232 => "0100000000000000",
  1233 => "0100000000000000",
  1234 => "0100000000000000",
  1235 => "0100000000000000",
  1236 => "0100000000000000",
  1237 => "0100000000000000",
  1238 => "0100000000000000",
  1239 => "0100000000000000",
  1240 => "0100000000000000",
  1241 => "0100000000000000",
  1242 => "0100000000000000",
  1243 => "0100000000000000",
  1244 => "0100000000000000",
  1245 => "0100000000000000",
  1246 => "0100000000000000",
  1247 => "0100000000000000",
  1248 => "0100000000000000",
  1249 => "0100000000000000",
  1250 => "0100000000000000",
  1251 => "0100000000000000",
  1252 => "0100000000000000",
  1253 => "0100000000000000",
  1254 => "0100000000000000",
  1255 => "0100000000000000",
  1256 => "0100000000000000",
  1257 => "0100000000000000",
  1258 => "0100000000000000",
  1259 => "0100000000000000",
  1260 => "0100000000000000",
  1261 => "0100000000000000",
  1262 => "0100000000000000",
  1263 => "0100000000000000",
  1264 => "0100000000000000",
  1265 => "0100000000000000",
  1266 => "0100000000000000",
  1267 => "0100000000000000",
  1268 => "0100000000000000",
  1269 => "0100000000000000",
  1270 => "0100000000000000",
  1271 => "0100000000000000",
  1272 => "0100000000000000",
  1273 => "0100000000000000",
  1274 => "0100000000000000",
  1275 => "0100000000000000",
  1276 => "0100000000000000",
  1277 => "0100000000000000",
  1278 => "0100000000000000",
  1279 => "0100000000000000",
  1280 => "0100000000000000",
  1281 => "0100000000000000",
  others => "0100000000000000"
  
  ); 
signal read_data_1,read_data_2,read_ins : std_logic_vector(15 downto 0);

begin
process(RAM_CLOCK)is
begin
 if(rising_edge(RAM_CLOCK)) then
    if(RAM_DATA_WR='1') then  
      RAM(to_integer(unsigned(RAM_DATA_ADDR))-1) <= RAM_DATA_IN(15 downto 0);
      RAM(to_integer(unsigned(RAM_DATA_ADDR))) <= RAM_DATA_IN(31 downto 16);
    end if;
    if(RAM_INS_WR='1') then  
      RAM(to_integer(unsigned(RAM_INS_ADDR))) <= RAM_INS_IN;
    end if;

 end if;  

end process;

read_data_2 <= RAM(to_integer(unsigned(RAM_DATA_ADDR))) when RAM_DATA_ADDR /= "UUUUUUUUUUU" else (others => 'Z');
-- ezzzzzaaaaat
read_data_1 <= RAM(to_integer(unsigned(RAM_DATA_ADDR)) - 1) when RAM_DATA_ADDR /= "UUUUUUUUUUU" and RAM_DATA_ADDR /= "00000000000" else (others => 'Z');

read_ins <=RAM(to_integer(unsigned(RAM_INS_ADDR))) when RAM_INS_ADDR /= "UUUUUUUUUUU" else "0100000000000000";

RAM_INS_OUT<=read_ins;
RAM_DATA_OUT<=read_data_2 & read_data_1;
end Behavioral;

